package ahb_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "ahb_agent_config.sv"
    `include "ahb_transaction.sv"
    `include "ahb_sequencer.sv"
    `include "ahb_driver.sv"
    `include "ahb_monitor.sv"
    `include "ahb_agent_active.sv"
    `include "ahb_monitor_passive.sv"
    `include "ahb_agent_passive.sv"
endpackage: ahb_pkg


package test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import ahb_pkg::*;
    import ahb_sequences_pkg::*;
    import apb_pkg::apb_sequence;
    import env_pkg::*;

    `include "ahb_apb_vseq.sv"
    `include "base_test.sv"
    `include "init_vseq_from_test.sv"

endpackage: test_pkg


package apb_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "apb_slave.sv"
    `include "apb_agent_config.sv"
    `include "apb_transaction.sv"
    `include "apb_sequencer.sv"
    `include "apb_sequence.sv"
    `include "apb_driver.sv"
    `include "apb_monitor.sv"
    `include "apb_agent.sv"
endpackage: apb_pkg

